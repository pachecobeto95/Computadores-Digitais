Entity FFJK_PR_CLR is port(j, k, clk, pr, clr : in bit;
                            q : out bit
                    );
End FFJK_PR_CLR;



Architecture Hybrid of FFJK_PR_CLR is 

Component FFJK
  port (j, k, clk : in bit;
                        q, nq : out bit
                );
End Component;

signal qt : bit;

Begin
  
  FFJK0 : FFJK port map(j, k, clk, qt);
  
  q <= '1' when (clr = '1') and (pr = '0') else
        '0' when (clr = '0') and (pr = '1') else
        qt;  
  
  
  
  
  
End Hybrid;
