Entity DETECTOR is port(x, clk : in bit;
                          z : out bit
                  );
End DETECTOR;



Architecture Comportamental of DETECTOR is
  Type estado is (reset, tem1, tem10, tem101, tem1011);
    
  signal atual : estado := reset;
  
  Begin
  
    Saida : Process(atual)
    
    Begin
      
        if (atual = tem1011) then z <= '1';
        else z <= '0';
        end if;   
    
    End Process;
    
    Transition : Process(clk)
    
    Begin
      
      if (clk'Event) and (clk = '1') then
        case atual is
        
          when reset => if (x = '1') then 
                          atual <= tem1;
                        end if;
                          
          when tem1 =>  if (x = '0') then
                          atual <= tem10;
                        end if;
                      
          when tem10 => if (x = '0') then
                          atual <= reset;
                        else 
                          atual <= tem101; 
                        end if;
                                 
          when tem101 => if (x = '0') then
                            atual <= tem10;
                         else
                            atual <= tem1011;
                         end if;
          when tem1011 => if (x = '0') then
                            atual <= tem10;
                          else 
                            atual <= tem1;
                          end if;               
       end case; 
      
        
      end if;
  
    End Process;
  
  
  
  
  
  End Comportamental;  
